module circuit2(
    input A,
    input B,
    output F
);
    and (F, A, B); // F = A AND B
endmodule
